package pack;
    `include "transaction.svh";
    `include "sequencer.svh";
    `include "driver.svh";
    `include "monitor.svh";
    `include "scoreboard.svh";
    `include "subscriber.svh";
    `include "environment.svh";
endpackage